----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:39:35 10/26/2018 
-- Design Name: 
-- Module Name:    prototip_1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity prototip_1 is
    Port ( iA : in  STD_LOGIC;
           iB : in  STD_LOGIC;
           iC : in  STD_LOGIC;
           oS : out  STD_LOGIC;
           oC : out  STD_LOGIC);
end prototip_1;

architecture Behavioral of prototip_1 is

begin

oS <= (iA xor iB) xor iC;
oC <= ((iA xor iB) and iC) or (iA and iB);

end Behavioral;

